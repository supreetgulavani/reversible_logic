/////////////////////////////////////////////////////////////////////
//  Filename: toffoli_gate.sv
//  
//  An Implementation of Toffoli Gate in SystemVerilog
//  
//  Author: Supreet Gulavani
//  05/22/2025
/////////////////////////////////////////////////////////////////////

module toffoli_gate(A, B, C, P, Q, R);

    input logic A;
    input logic B;
    input logic C;
    output logic P;
    output logic Q;
    output logic R;

    assign P = A;
    assign Q = B;
    assign R = (A & B) ^ C;

endmodule